library verilog;
use verilog.vl_types.all;
entity fmat_alu_testbench is
end fmat_alu_testbench;
