library verilog;
use verilog.vl_types.all;
entity fetchUnit_testbench is
end fetchUnit_testbench;
