module to_flag (
	input [7:0] input_i,
	output output_o);
	
assign output_o = input_i[0];

endmodule