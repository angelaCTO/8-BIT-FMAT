library verilog;
use verilog.vl_types.all;
entity p3_testbench is
end p3_testbench;
