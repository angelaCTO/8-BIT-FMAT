module p3_testbench();
// Declare inputs as regs and outputs as wires

	reg clk;			        // Clock 
	reg start_i;            // flag: whether to jump to the start address
	reg [7:0] start_addr_i; // the address of the beginning of the program
	wire writeEnable_o;
	wire [3:0] regWrite_o;
	wire [7:0] dataWrite_o;
	wire [7:0] instr_o;
	wire [7:0] pc_o;
	wire halt_o;
	wire yesJump_o;
	wire [7:0] target_o;
	
// Initialize all variables
initial begin        
	clk = 1;       // initial value of clock
	start_i = 0;
	start_addr_i = 0;
	
	
	#10 start_i = 1;
	#10 start_i = 0;
end

 // Clock generator
always begin
   #5  clk = ~clk; // Toggle clock every 5 ticks
						// this makes the clock cycle 10 ticks
end

// the following creates an instance of our program_counter register.
//   I copied this code verbatim from the walkthough.v that was
//   generated by Quartus when I created the .v file from the .bdf.

p2 b2v_inst(
	.clk(clk),
	.start_i(start_i),
	.start_addr_i(start_addr_i),
	.writeEnable_o(writeEnable_o),
	.regWrite_o(regWrite_o),
	.dataWrite_o(dataWrite_o),
	.instr_o(instr_o),
	.pc_o(pc_o),
	.halt_o(halt_o),
	.yesJump_o(yesJump_o),
	.target_o(target_o)
);
endmodule
